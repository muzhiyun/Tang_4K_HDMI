//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.09 Education
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Sun Apr 23 16:46:39 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [2:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [1:1] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [2:2] prom_inst_2_dout;
wire [28:0] prom_inst_3_dout_w;
wire [2:0] prom_inst_3_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_1.INIT = 16'h0200;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFC00000000FFFFFFFC0000000000000000FFFFFFFC00000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h00000000000000000000FFFFFFFC00000000000000000000000000000000FFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000FFFFFFFC00000000000000000000000000000000FFFFFFFC000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000FFFFFFFC0000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h000000000000FFFFFFFC00000000000000000000000000000000FFFFFFFC0000;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFC00000000000000000000000000000000FFFFFFFC00000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h000000000000000000000000000400000000000000000000000000000000FFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFE0000000000000000000001E0000000007FFFFFFE0000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h000000000000000003000FFFFFFFE0000000000000000000000FFFFFFF800FFF;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000FFFFFFFE00000000000000000000000000001000FFFFFFFE00000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000000000000000000000000FFFFFFFE000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000FFFFFFFE00000000000000000000000000000000FFFFFFFE000;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFE00000000000000000000000000000000FFFFFFFE0000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h000000000000000000000FFFFFFFE00000000000000000000000000000000FFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFC0000000000000000000000000000000000000FF80000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h00000000000000000000000001EFFC4400000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h000003FFF0000000000000000000000000000000000000007000000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'hFF003E1F01F8000030F90E000000038F00E00001F000083801F00000007E1F00;
defparam prom_inst_0.INIT_RAM_29 = 256'hE03C1E000000010780E3C01FFF807F9E031803FFE0FCCE000000010700E3F007;
defparam prom_inst_0.INIT_RAM_2A = 256'h80E0E07FFFE0385E070C0780F0003E000000000780E1C03FFFC07C4E020807EB;
defparam prom_inst_0.INIT_RAM_2B = 256'h0F0400FEF01E3C0000000FE7C0F0F07FFFE0007E07FC0383F003FE00000003C7;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000070780F078FFFFF03E1C0E02001E707C1C0000000787807070FFFFF00FFE;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFE0F83F3E038FBC707C3D000000019E00FC787FFFE0781C0E010F1C70783F00;
defparam prom_inst_0.INIT_RAM_2E = 256'hDC000000000000000010F03FFFE07C3800080E3CF80000000000000001F2F87F;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000FFF0000000000000000000000000000000000003FFFE00000000003F8;
defparam prom_inst_0.INIT_RAM_30 = 256'h00000000000000000000000000000003FC000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000003C00000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h00000000FF80000000000000000000000000000000000000FF00000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h00000000000000000000000000000001FFC00000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000FF80000000000000000000000000000000000001FFC00000;
defparam prom_inst_0.INIT_RAM_3C = 256'h3C00000000000000000000000000000000000000FF0000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFF000000000FFFFFFFC0000000000000000FFFFFFFC00000000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFC00000000000000000000000000000000FFFFFFFC00000000000000001FFF;
defparam prom_inst_1.INIT_RAM_0D = 256'h00000000000000000000FFFFFFFC00000000000000000000000000000000FFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'h0000FFFFFFFC00000000000000000000000000000000FFFFFFFC000000000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000BFFFFFFC0000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_10 = 256'h000000000000FFFFFFFC00000000000000000000000000000000FFFFFFFC0000;
defparam prom_inst_1.INIT_RAM_11 = 256'h001400000000000000000000000000000000E1E71E9C00000000000000000000;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFE0000000000000000000001FFFFFFF0007FFFFFFC0000000000000000000;
defparam prom_inst_1.INIT_RAM_13 = 256'h00000000001FFFFFFF800FFFFFFFE0000000000000000000001FFFFFFF800FFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFF800FFFFFFFE0000000000000000000001FFFFFFF800FFFFFFFE00000000000;
defparam prom_inst_1.INIT_RAM_15 = 256'h0000000000000000001FFFFFFF800FFFFFFFE0000000000000000000001FFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'h001FFFFFFF800FFFFFFFE0000000000000000000001FFFFFFF800FFFFFFFE000;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFE0000000000000000000001FFFFFFF800FFFFFFFE0000000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h00000000001FFFFFFF800FFFFFFFE0000000000000000000001FFFFFFF800FFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFC00000000000000000000000000000001FF801FF80000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h000000000000000000000001FFFFFFFC00000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_1B = 256'h00000001FFFFFFFC00000000000000000000000000000001FFFFFFFC00000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h00000000000000000000000000000001FFFFFFFC000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000001FFFFFFFC00000000000000000000000000000001FFFFFFFC;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFC00000000000000000000000000000001FFFFFFFC0000000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h000000000000000000000001FFFFFFFC00000000000000000000000000000001;
defparam prom_inst_1.INIT_RAM_20 = 256'h000000000000000000000000000000000000000000000001FFFFFFFC00000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h000003FFF0000000000000000000000000000000000000007000000000000000;
defparam prom_inst_1.INIT_RAM_28 = 256'hFF003E1F01F8000030F90E000000038F00E00001F000083801F00000007E1F00;
defparam prom_inst_1.INIT_RAM_29 = 256'hE03C1E000000010780E3C01FFF807F9E031803FFE0FCCE000000010700E3F007;
defparam prom_inst_1.INIT_RAM_2A = 256'h80E0E07FFFE0385E070C0780F0003E000000000780E1C03FFFC07C4E020807EB;
defparam prom_inst_1.INIT_RAM_2B = 256'h0F0400FEF01E3C0000000FE7C0F0F07FFFE0007E07FC0383F003FE00000003C7;
defparam prom_inst_1.INIT_RAM_2C = 256'h0000070780F078FFFFF03E1C0E02001E707C1C0000000787807070FFFFF00FFE;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFE0F83F3E038FBC707C3D000000019E00FC787FFFE0781C0E010F1C70783F00;
defparam prom_inst_1.INIT_RAM_2E = 256'hDC000000000000000010F03FFFE07C3800080E3CF80000000000000001F2F87F;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000FFF0000000000000000000000000000000000003FFFE00000000003F8;
defparam prom_inst_1.INIT_RAM_30 = 256'h00000000000000000000000000000003FC000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000003C00000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h00000000FF80000000000000000000000000000000000000FF00000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h00000000000000000000000000000001FFC00000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000FF80000000000000000000000000000000000001FFC00000;
defparam prom_inst_1.INIT_RAM_3C = 256'h3C00000000000000000000000000000000000000FF0000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFC00000000FFFFFFFC0000000000000000FFFFFFFC00000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFC0000000000000000FFFFFFFC00000001FFFFFFFC0000000000000000FFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'h0000FFFFFFFC00000001FFFFFFFC0000000000000001FFFFFFFC00000001FFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'h0001FFFFFFFC0000000000000001FFFFFFFC00000001FFFFFFFC000000000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h000000000000FFFFFFFC00000001FFFFFFFC0000000000000000FFFFFFFC0000;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFC00000001FFFFFFFC0000000000000000FFFFFFFC00000001FFFFFFFC0000;
defparam prom_inst_2.INIT_RAM_11 = 256'h003C00000000000000000000000400000001FFFFFFFC0000000000000000FFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFE0000000000000000000001E0000000000000003E0000000000000002000;
defparam prom_inst_2.INIT_RAM_13 = 256'h000000000000000000000FFFFFFFE0000000000000000000000FFFFFFF800FFF;
defparam prom_inst_2.INIT_RAM_14 = 256'h00000FFFFFFFE00000000000000000000000000000000FFFFFFFE00000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h00000000000000000000000000000FFFFFFFE000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0000000000000FFFFFFFE00000000000000000000000000000000FFFFFFFE000;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFE00000000000000000000000000000000FFFFFFFE0000000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h000000000000000000000FFFFFFFE00000000000000000000000000000000FFF;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFFFFC0000000000000000000000000000000000801FF80000000000000000;
defparam prom_inst_2.INIT_RAM_1A = 256'h000000000000000000000000FFFFFFFC00000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_1B = 256'h00000001FFFFFFFC00000000000000000000000000000001FFFFFFFC00000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h00000000000000000000000000000001FFFFFFFC000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0000000000000001FFFFFFFC00000000000000000000000000000001FFFFFFFC;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFFFFC00000000000000000000000000000001FFFFFFFC0000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h000000000000000000000001FFFFFFFC00000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_20 = 256'h000000000000000000000000000000000000000000000001FFFFFFFC00000000;
defparam prom_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_27 = 256'h000003FFF0000000000000000000000000000000000000007000000000000000;
defparam prom_inst_2.INIT_RAM_28 = 256'hFF003E1F01F8000030F90E000000038F00E00001F000083801F00000007E1F00;
defparam prom_inst_2.INIT_RAM_29 = 256'hE03C1E000000010780E3C01FFF807F9E031803FFE0FCCE000000010700E3F007;
defparam prom_inst_2.INIT_RAM_2A = 256'h80E0E07FFFE0385E070C0780F0003E000000000780E1C03FFFC07C4E020807EB;
defparam prom_inst_2.INIT_RAM_2B = 256'h0F0400FEF01E3C0000000FE7C0F0F07FFFE0007E07FC0383F003FE00000003C7;
defparam prom_inst_2.INIT_RAM_2C = 256'h0000070780F078FFFFF03E1C0E02001E707C1C0000000787807070FFFFF00FFE;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFE0F83F3E038FBC707C3D000000019E00FC787FFFE0781C0E010F1C70783F00;
defparam prom_inst_2.INIT_RAM_2E = 256'hDC000000000000000010F03FFFE07C3800080E3CF80000000000000001F2F87F;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000FFF0000000000000000000000000000000000003FFFE00000000003F8;
defparam prom_inst_2.INIT_RAM_30 = 256'h00000000000000000000000000000003FC000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000001800000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h00000000FF800000000000000000000000000000000000007F00000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h00000000000000000000000000000001FF800000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000FF80000000000000000000000000000000000001FF800000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000FF0000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[28:0],prom_inst_3_dout[2:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 4;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h4444444444444444444444444444440000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000004;
defparam prom_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000444444444444444444444444444444400;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_4 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(dout[1]),
  .I0(prom_inst_1_dout[1]),
  .I1(prom_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[2]),
  .I0(prom_inst_2_dout[2]),
  .I1(prom_inst_3_dout[2]),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM
